library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity BinDecROM is
    port(
        reset : in std_logic;
        address : in std_logic_vector(7 downto 0);
                                                
        dataOut : out std_logic_vector(7 downto 0)
    );
end BinDecROM;

architecture behavioral of BinDecROM is 
type rom_type is array (0 to 255) of std_logic_vector(7 downto 0);
signal BinDecROM : rom_type := (
    X"00",
    X"01",
    X"02",
    X"03",
    X"04",
    X"05",
    X"06",
    X"07",
    X"08",
    X"09",
    X"10",
    X"11",
    X"12",
    X"13",
    X"14",
    X"15",
    X"16",
    X"17",
    X"18",
    X"19",
    X"20",
    X"21",
    X"22",
    X"23",
    X"24",
    X"25",
    X"26",
    X"27",
    X"28",
    X"29",
    X"30",
    X"31",
    X"32",
    X"33",
    X"34",
    X"35",
    X"36",
    X"37",
    X"38",
    X"39",
    X"40",
    X"41",
    X"42",
    X"43",
    X"44",
    X"45",
    X"46",
    X"47",
    X"48",
    X"49",
    X"50",
    X"51",
    X"52",
    X"53",
    X"54",
    X"55",
    X"56",
    X"57",
    X"58",
    X"59",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00",
    X"00"
);

--attribute rom_style : string;
--attribute rom_style of BinDecROM : signal is "block";-- block dice al tool di sintesi di inferire blocchi di RAMB, 
--                                               -- distributed di usare le LUT
begin

process(address)
  begin
    if (reset = '1') then
       dataOut <= BinDecROM(conv_integer("00000000"));
    else
        dataOut <= BinDecROM(conv_integer(address));
    end if;
    
end process;
end behavioral;