library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity EncoderDecimalBCD is
    port(
        input: in std_logic_vector(0 to 5);
        
        output: out std_logic_vector(7 downto 0)
    );
end EncoderDecimalBCD;

architecture Dataflow of EncoderDecimalBCD is

begin
    with input select
        output <=   "00000000" when "000000",
                    "00000001" when "000001",
                    "00000010" when "000010",
                    "00000011" when "000011",
                    "00000100" when "000100",
                    "00000101" when "000101",
                    "00000110" when "000110",
                    "00000111" when "000111",
                    "00001000" when "001000",
                    "00001001" when "001001",
                    "00010000" when "001010",
                    "00010001" when "001011",
                    "00010010" when "001100",
                    "00010011" when "001101",
                    "00010100" when "001110",
                    "00010101" when "001111",
                    "00010110" when "010000",
                    "00010111" when "010001",
                    "00011000" when "010010",
                    "00011001" when "010011",
                    "00100000" when "010100",
                    "00100001" when "010101",
                    "00100010" when "010110",
                    "00100011" when "010111",
                    "00100100" when "011000",
                    "00100101" when "011001",
                    "00100110" when "011010",
                    "00100111" when "011011",
                    "00101000" when "011100",
                    "00101001" when "011101",
                    "00110000" when "011110",
                    "00110001" when "011111",
                    "00110010" when "100000",
                    "00110011" when "100001",
                    "00110100" when "100010",
                    "00110101" when "100011",
                    "00110110" when "100100",
                    "00110111" when "100101",
                    "00111000" when "100110",
                    "00111001" when "100111",
                    "01000000" when "101000",
                    "01000001" when "101001",
                    "01000010" when "101010",
                    "01000011" when "101011",
                    "01000100" when "101100",
                    "01000101" when "101101",
                    "01000110" when "101110",
                    "01000111" when "101111",
                    "01001000" when "110000",
                    "01001001" when "110001",
                    "01010000" when "110010",
                    "01010001" when "110011",
                    "01010010" when "110100",
                    "01010011" when "110101",
                    "01010100" when "110110",
                    "01010101" when "110111",
                    "01010110" when "111000",
                    "01010111" when "111001",
                    "01011000" when "111010",
                    "01011001" when "111011",
                    "01100000" when "111100",
                    "01100001" when "111101",
                    "01100010" when "111110",
                    "01100011" when "111111",
                    "11111111" when others;

end Dataflow;
