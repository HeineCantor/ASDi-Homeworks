library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity EncoderSignedBCD is
    port(
        input: in std_logic_vector(7 downto 0);
        
        output: out std_logic_vector(15 downto 0)
    );
end EncoderSignedBCD;

architecture Dataflow of EncoderSignedBCD is

begin
    with input select
        output <=   "0000000000000000" when "00000000",
                    "0000000000000001" when "00000001",
                    "0000000000000010" when "00000010",
                    "0000000000000011" when "00000011",
                    "0000000000000100" when "00000100",
                    "0000000000000101" when "00000101",
                    "0000000000000110" when "00000110",
                    "0000000000000111" when "00000111",
                    "0000000000001000" when "00001000",
                    "0000000000001001" when "00001001",
                    "0000000000010000" when "00001010",
                    "0000000000010001" when "00001011",
                    "0000000000010010" when "00001100",
                    "0000000000010011" when "00001101",
                    "0000000000010100" when "00001110",
                    "0000000000010101" when "00001111",
                    "0000000000010110" when "00010000",
                    "0000000000010111" when "00010001",
                    "0000000000011000" when "00010010",
                    "0000000000011001" when "00010011",
                    "0000000000100000" when "00010100",
                    "0000000000100001" when "00010101",
                    "0000000000100010" when "00010110",
                    "0000000000100011" when "00010111",
                    "0000000000100100" when "00011000",
                    "0000000000100101" when "00011001",
                    "0000000000100110" when "00011010",
                    "0000000000100111" when "00011011",
                    "0000000000101000" when "00011100",
                    "0000000000101001" when "00011101",
                    "0000000000110000" when "00011110",
                    "0000000000110001" when "00011111",
                    "0000000000110010" when "00100000",
                    "0000000000110011" when "00100001",
                    "0000000000110100" when "00100010",
                    "0000000000110101" when "00100011",
                    "0000000000110110" when "00100100",
                    "0000000000110111" when "00100101",
                    "0000000000111000" when "00100110",
                    "0000000000111001" when "00100111",
                    "0000000001000000" when "00101000",
                    "0000000001000001" when "00101001",
                    "0000000001000010" when "00101010",
                    "0000000001000011" when "00101011",
                    "0000000001000100" when "00101100",
                    "0000000001000101" when "00101101",
                    "0000000001000110" when "00101110",
                    "0000000001000111" when "00101111",
                    "0000000001001000" when "00110000",
                    "0000000001001001" when "00110001",
                    "0000000001010000" when "00110010",
                    "0000000001010001" when "00110011",
                    "0000000001010010" when "00110100",
                    "0000000001010011" when "00110101",
                    "0000000001010100" when "00110110",
                    "0000000001010101" when "00110111",
                    "0000000001010110" when "00111000",
                    "0000000001010111" when "00111001",
                    "0000000001011000" when "00111010",
                    "0000000001011001" when "00111011",
                    "0000000001100000" when "00111100",
                    "0000000001100001" when "00111101",
                    "0000000001100010" when "00111110",
                    "0000000001100011" when "00111111",
                    "0000000001100100" when "01000000",
                    "0000000001100101" when "01000001",
                    "0000000001100110" when "01000010",
                    "0000000001100111" when "01000011",
                    "0000000001101000" when "01000100",
                    "0000000001101001" when "01000101",
                    "0000000001110000" when "01000110",
                    "0000000001110001" when "01000111",
                    "0000000001110010" when "01001000",
                    "0000000001110011" when "01001001",
                    "0000000001110100" when "01001010",
                    "0000000001110101" when "01001011",
                    "0000000001110110" when "01001100",
                    "0000000001110111" when "01001101",
                    "0000000001111000" when "01001110",
                    "0000000001111001" when "01001111",
                    "0000000010000000" when "01010000",
                    "0000000010000001" when "01010001",
                    "0000000010000010" when "01010010",
                    "0000000010000011" when "01010011",
                    "0000000010000100" when "01010100",
                    "0000000010000101" when "01010101",
                    "0000000010000110" when "01010110",
                    "0000000010000111" when "01010111",
                    "0000000010001000" when "01011000",
                    "0000000010001001" when "01011001",
                    "0000000010010000" when "01011010",
                    "0000000010010001" when "01011011",
                    "0000000010010010" when "01011100",
                    "0000000010010011" when "01011101",
                    "0000000010010100" when "01011110",
                    "0000000010010101" when "01011111",
                    "0000000010010110" when "01100000",
                    "0000000010010111" when "01100001",
                    "0000000010011000" when "01100010",
                    "0000000010011001" when "01100011",
                    "0000000100000000" when "01100100",
                    "0000000100000001" when "01100101",
                    "0000000100000010" when "01100110",
                    "0000000100000011" when "01100111",
                    "0000000100000100" when "01101000",
                    "0000000100000101" when "01101001",
                    "0000000100000110" when "01101010",
                    "0000000100000111" when "01101011",
                    "0000000100001000" when "01101100",
                    "0000000100001001" when "01101101",
                    "0000000100010000" when "01101110",
                    "0000000100010001" when "01101111",
                    "0000000100010010" when "01110000",
                    "0000000100010011" when "01110001",
                    "0000000100010100" when "01110010",
                    "0000000100010101" when "01110011",
                    "0000000100010110" when "01110100",
                    "0000000100010111" when "01110101",
                    "0000000100011000" when "01110110",
                    "0000000100011001" when "01110111",
                    "0000000100100000" when "01111000",
                    "0000000100100001" when "01111001",
                    "0000000100100010" when "01111010",
                    "0000000100100011" when "01111011",
                    "0000000100100100" when "01111100",
                    "0000000100100101" when "01111101",
                    "0000000100100110" when "01111110",
                    "0000000100100111" when "01111111",
                    "1111000100101000" when "10000000",
                    "1111000100100111" when "10000001",
                    "1111000100100110" when "10000010",
                    "1111000100100101" when "10000011",
                    "1111000100100100" when "10000100",
                    "1111000100100011" when "10000101",
                    "1111000100100010" when "10000110",
                    "1111000100100001" when "10000111",
                    "1111000100100000" when "10001000",
                    "1111000100011001" when "10001001",
                    "1111000100011000" when "10001010",
                    "1111000100010111" when "10001011",
                    "1111000100010110" when "10001100",
                    "1111000100010101" when "10001101",
                    "1111000100010100" when "10001110",
                    "1111000100010011" when "10001111",
                    "1111000100010010" when "10010000",
                    "1111000100010001" when "10010001",
                    "1111000100010000" when "10010010",
                    "1111000100001001" when "10010011",
                    "1111000100001000" when "10010100",
                    "1111000100000111" when "10010101",
                    "1111000100000110" when "10010110",
                    "1111000100000101" when "10010111",
                    "1111000100000100" when "10011000",
                    "1111000100000011" when "10011001",
                    "1111000100000010" when "10011010",
                    "1111000100000001" when "10011011",
                    "1111000100000000" when "10011100",
                    "1111000010011001" when "10011101",
                    "1111000010011000" when "10011110",
                    "1111000010010111" when "10011111",
                    "1111000010010110" when "10100000",
                    "1111000010010101" when "10100001",
                    "1111000010010100" when "10100010",
                    "1111000010010011" when "10100011",
                    "1111000010010010" when "10100100",
                    "1111000010010001" when "10100101",
                    "1111000010010000" when "10100110",
                    "1111000010001001" when "10100111",
                    "1111000010001000" when "10101000",
                    "1111000010000111" when "10101001",
                    "1111000010000110" when "10101010",
                    "1111000010000101" when "10101011",
                    "1111000010000100" when "10101100",
                    "1111000010000011" when "10101101",
                    "1111000010000010" when "10101110",
                    "1111000010000001" when "10101111",
                    "1111000010000000" when "10110000",
                    "1111000001111001" when "10110001",
                    "1111000001111000" when "10110010",
                    "1111000001110111" when "10110011",
                    "1111000001110110" when "10110100",
                    "1111000001110101" when "10110101",
                    "1111000001110100" when "10110110",
                    "1111000001110011" when "10110111",
                    "1111000001110010" when "10111000",
                    "1111000001110001" when "10111001",
                    "1111000001110000" when "10111010",
                    "1111000001101001" when "10111011",
                    "1111000001101000" when "10111100",
                    "1111000001100111" when "10111101",
                    "1111000001100110" when "10111110",
                    "1111000001100101" when "10111111",
                    "1111000001100100" when "11000000",
                    "1111000001100011" when "11000001",
                    "1111000001100010" when "11000010",
                    "1111000001100001" when "11000011",
                    "1111000001100000" when "11000100",
                    "1111000001011001" when "11000101",
                    "1111000001011000" when "11000110",
                    "1111000001010111" when "11000111",
                    "1111000001010110" when "11001000",
                    "1111000001010101" when "11001001",
                    "1111000001010100" when "11001010",
                    "1111000001010011" when "11001011",
                    "1111000001010010" when "11001100",
                    "1111000001010001" when "11001101",
                    "1111000001010000" when "11001110",
                    "1111000001001001" when "11001111",
                    "1111000001001000" when "11010000",
                    "1111000001000111" when "11010001",
                    "1111000001000110" when "11010010",
                    "1111000001000101" when "11010011",
                    "1111000001000100" when "11010100",
                    "1111000001000011" when "11010101",
                    "1111000001000010" when "11010110",
                    "1111000001000001" when "11010111",
                    "1111000001000000" when "11011000",
                    "1111000000111001" when "11011001",
                    "1111000000111000" when "11011010",
                    "1111000000110111" when "11011011",
                    "1111000000110110" when "11011100",
                    "1111000000110101" when "11011101",
                    "1111000000110100" when "11011110",
                    "1111000000110011" when "11011111",
                    "1111000000110010" when "11100000",
                    "1111000000110001" when "11100001",
                    "1111000000110000" when "11100010",
                    "1111000000101001" when "11100011",
                    "1111000000101000" when "11100100",
                    "1111000000100111" when "11100101",
                    "1111000000100110" when "11100110",
                    "1111000000100101" when "11100111",
                    "1111000000100100" when "11101000",
                    "1111000000100011" when "11101001",
                    "1111000000100010" when "11101010",
                    "1111000000100001" when "11101011",
                    "1111000000100000" when "11101100",
                    "1111000000011001" when "11101101",
                    "1111000000011000" when "11101110",
                    "1111000000010111" when "11101111",
                    "1111000000010110" when "11110000",
                    "1111000000010101" when "11110001",
                    "1111000000010100" when "11110010",
                    "1111000000010011" when "11110011",
                    "1111000000010010" when "11110100",
                    "1111000000010001" when "11110101",
                    "1111000000010000" when "11110110",
                    "1111000000001001" when "11110111",
                    "1111000000001000" when "11111000",
                    "1111000000000111" when "11111001",
                    "1111000000000110" when "11111010",
                    "1111000000000101" when "11111011",
                    "1111000000000100" when "11111100",
                    "1111000000000011" when "11111101",
                    "1111000000000010" when "11111110",
                    "1111000000000001" when "11111111",
                    "11111111" when others;

end Dataflow;
